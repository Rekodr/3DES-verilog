`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/06/2019 04:53:14 PM
// Design Name: 
// Module Name: round_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module round_tb();

reg clk;
reg [31:0] R0;
wire [31:0] R1;
wire [31:0] R2;
wire [31:0] R3;
wire [31:0] R4;
wire [31:0] R5;
wire [31:0] R6;
wire [31:0] R7;
wire [31:0] R8;
wire [31:0] R9;
wire [31:0] R10;
wire [31:0] R11;
wire [31:0] R12;
wire [31:0] R13;
wire [31:0] R14;
wire [31:0] R15;
wire [31:0] R16;

reg [31:0] L0;
wire [31:0] L1;
wire [31:0] L2;
wire [31:0] L3;
wire [31:0] L4;
wire [31:0] L5;
wire [31:0] L6;
wire [31:0] L7;
wire [31:0] L8;
wire [31:0] L9;
wire [31:0] L10;
wire [31:0] L11;
wire [31:0] L12;
wire [31:0] L13;
wire [31:0] L14;
wire [31:0] L15;
wire [31:0] L16;


reg [47:0] K1;
reg [47:0] K2;
reg [47:0] K3;
reg [47:0] K4;
reg [47:0] K5;
reg [47:0] K6;
reg [47:0] K7;
reg [47:0] K8;
reg [47:0] K9;
reg [47:0] K10;
reg [47:0] K11;
reg [47:0] K12;
reg [47:0] K13;
reg [47:0] K14;
reg [47:0] K15;
reg [47:0] K16;

round Rnd1(clk, L0, R0, K1, 1'b1, L1, R1);
round Rnd2(clk, L1, R1, K2, 1'b1, L2, R2);
round Rnd3(clk, L2, R2, K3, 1'b1, L3, R3);
round Rnd4(clk, L3, R3, K4, 1'b1, L4, R4);
round Rnd5(clk, L4, R4, K5, 1'b1, L5, R5);
round Rnd6(clk, L5, R5, K6, 1'b1, L6, R6);
round Rnd7(clk, L6, R6, K7, 1'b1, L7, R7);
round Rnd8(clk, L7, R7, K8, 1'b1, L8, R8);
round Rnd9(clk, L8, R8, K9, 1'b1, L9, R9);
round Rnd10(clk, L9, R9, K10, 1'b1, L10, R10);
round Rnd11(clk, L10, R10, K11, 1'b1, L11, R11);
round Rnd12(clk, L11, R11, K12, 1'b1, L12, R12);
round Rnd13(clk, L12, R12, K13, 1'b1, L13, R13);
round Rnd14(clk, L13, R13, K14, 1'b1, L14, R14);
round Rnd15(clk, L14, R14, K15, 1'b1, L15, R15);
round Rnd16(clk, L15, R15, K16, 1'b0, L16, R16);

always #10 clk = ~clk;

initial 
begin
    clk = 0;
    K1 = 48'b000110_110000_001011_101111_111111_000111_000001_110010;
    K2 = 48'b011110_011010_111011_011001_110110_111100_100111_100101;
    K3 = 48'b010101_011111_110010_001010_010000_101100_111110_011001;
    K4 = 48'b011100_101010_110111_010110_110110_110011_010100_011101;
    K5 = 48'b011111_001110_110000_000111_111010_110101_001110_101000;
    K6 = 48'b011000_111010_010100_111110_010100_000111_101100_101111;
    K7 = 48'b111011_001000_010010_110111_111101_100001_100010_111100;
    K8 = 48'b111101_111000_101000_111010_110000_010011_101111_111011;
    K9 = 48'b111000_001101_101111_101011_111011_011110_011110_000001;
    K10 = 48'b101100_011111_001101_000111_101110_100100_011001_001111;
    K11 = 48'b001000_010101_111111_010011_110111_101101_001110_000110;
    K12 = 48'b011101_010111_000111_110101_100101_000110_011111_101001;
    K13 = 48'b100101_111100_010111_010001_111110_101011_101001_000001;
    K14 = 48'b010111_110100_001110_110111_111100_101110_011100_111010;
    K15 = 48'b101111_111001_000110_001101_001111_010011_111100_001010;
    K16 = 48'b110010_110011_110110_001011_000011_100001_011111_110101;
    
    #20;
    R0 = 32'b1111_0000_1010_1010_1111_0000_1010_1010;
    L0 = 32'b1100_1100_0000_0000_1100_1100_1111_1111;

end

endmodule
